module clockDivider(

input clk_in;
input clk_out;
);




if


//by default: period is 1 sec (1 HZ),
//have method to make it faster or slower
//can be either 1 HZ, 0.5 HZ (2 second period), 2 HZ (0.5 second period)