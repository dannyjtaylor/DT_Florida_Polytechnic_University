//Binary to Hex

module BinaryToHex(

input [3:0] bit1, bit2,
output 



endmodule

module convert(num);


	assign num = 1h'0 ? 8b'00000011 :
					 1h'1 ? 8b'10011111 :
					 1h'2 ? 8b'00100111 :
					 1h'3 ? 8b'00001101 :
					 1h'4 ? 8b'10011001 :
					 1h'5 ? 8b'01001101 :
					 1h'6 ? 8b'01000001 :
					 1h'7 ? 8b'00011111 :
					 1h'8 ? 8b'00000001 :
					 1h'9 ? 8b'00011001 :
	//				 1h'a ? 8b'
endmodule