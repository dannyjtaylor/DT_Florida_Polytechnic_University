/*module Add(input [3:0] A, B, output [3:0] sum);
	assign sum = A + B;
endmodule

module Multiply(input[3:0] A, B, output [7:0] product);
	assign product = A * B;
endmodule*/