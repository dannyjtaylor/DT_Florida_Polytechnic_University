module ShiftAndCombinehandson(

//FOR FPGA BOARD DATA DIRECTION
	//////////// SEG7 //////////
	output		     [7:0]		HEX0,
	output		     [7:0]		HEX1,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW);

endmodule
	